module datamem();


endmodule