module datamem();


endmodule
